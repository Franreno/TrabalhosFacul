*
v1 i 0 dc 6
r1 i 1 27k
r2 1 0 47k
*

.tran