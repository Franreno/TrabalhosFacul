Circuito Balun LC

Vin 1 0 AC 12 SIN(0 12 1024 0 0 90)


Rout 2 3 1483

L1 1 2 6.95436m
L2 3 0 6.95436m

C1 2 0 3.473u
C2 1 3 3.473u

.AC LIN 1 1024 1024
.print AC V(2) V(3)

.tran 1 20ms 10ms
.end







