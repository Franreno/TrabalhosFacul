Cir

v1 1 0 dc 0 ac 5

r1 1 2 200

l1 2 3 125m

c1 3 0 1u

.ac dec 10 1 1MEG

.print ac vdb(vout)
.plot ac vdb(vout)

.end