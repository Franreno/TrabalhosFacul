*Netlist do circuito. Trabalho SPICE-SEL0602. Francisco Reis Nogueira 11954374

V1 1 0 ac 7 SIN(0 7 47.1098631552 0 0 0)

r1 1 2 8

c1 2 3 0.04

r2 3 0 74

c2 3 4 0.02

r3 4 0 37

r4 4 5 5

l1 5 0 0.5

.AC LIN 1 47.11 47.11
.TRAN 1 12 10

.print AC V(3,0) VP(3,0) V(4,0) VP(4,0);
.print AC I(r2) IP(r2) I(r3) IP(r3) I(r4) IP(r4);

.probe

.end     