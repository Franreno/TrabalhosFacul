EXEMPLO 2 RESOLUCAO

V1 1 0 DC 24
R1 1 2 5
L1 2 3 1
C1 3 0 0.25

.IC I(L1) = 4
.IC v(3,0) = 4

.tran 0.05 1 uic
.plot tran I(R1)
.end