chave
*
v1 i 0 dc 24
r1 i o 6
r2 o 0 3
c1 o 0 2
*

*
.ic v(o) = 20
.ic i(o) = 0
*

*
.tran .1 20
*

.end
