EXEMPLO

V1 1 0 DC 100
R1 1 2 20
R2 2 0 30

.DC V1 100 100 1

.PRINT DC I(R1)
.PRINT DC V(1,2) V(2,0)

.END
